-----------------------------------------------------------
-- Entity Name: rtg_mux2to1_w4
-----------------------------------------------------------

library IEEE;
use IEEE.std_logic_1164.all;

entity rtg_mux2to1_w4 is
  port (
    SEL : in std_logic;
    DIN0 : in std_logic_vector(3 downto 0);
    DIN1 : in std_logic_vector(3 downto 0);
    DOUT : out std_logic_vector(3 downto 0)
  );
end entity rtg_mux2to1_w4;

architecture RTL of rtg_mux2to1_w4 is


begin
  DOUT <= DIN0 when SEL = '0' else 
	DIN1 when SEL = '1' else 
	"XXXX";
end RTL;

-----------------------------------------
-- Generated by ASIP Meister ver.1.1 --
-----------------------------------------
