-- VHDL       : '87
-- Module     : Sign Extender
-- Feature    : extend sign
-- References : Started from scratch.
-- Author     : Tak. Tokihisa
-- Version : 1.0  : 2002/01/14

-- Functionality : behavior level
--  port
--   data_in  : data extended
--   data_out : extended data 
--   mode     : 0  zero extention
--            : 1  sign extention

library IEEE;
  use IEEE.std_logic_1164.all;
  use IEEE.std_logic_unsigned.all;

entity fhm_extender_w28 is
  port (data_in  : in std_logic_vector(27 downto 0);
        mode     : in std_logic;
        data_out : out std_logic_vector(31 downto 0));
end fhm_extender_w28;

architecture behavior of fhm_extender_w28 is
begin
  process (data_in, mode)
    begin
      data_out(27 downto 0) <= data_in(27 downto 0);
      if mode = '0' then
        data_out(31 downto 28) <= "0000";
      else
        for i in 31 downto 28 loop
          data_out(i) <= data_in(27);
        end loop;
      end if;
  end process;
end behavior;

-----------------------------------------
-- Generated by ASIP Meister ver.1.1 --
-----------------------------------------
