library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.ALL;
use work.debounce_pack.ALL;
--fpga4student.com: FPGA projects, Verilog projects, VHDL projects
-- VHDL code for button debouncing on FPGA 
-- Testbench VHDL code for button debouncing
ENTITY tb_debouncer2 IS
END tb_debouncer2;
 
ARCHITECTURE behavior OF tb_debouncer2 IS
    -- Component Declaration for VHDL code for button debouncing
    COMPONENT debouncer2
    PORT(
         pbutton : IN  std_logic;
         clk : IN  std_logic;
--         rst : IN  std_logic;
         pd_deb : OUT  std_logic
        );
    END COMPONENT;
   signal pbutton : std_logic := '0';
   signal clk : std_logic := '0';
--   signal rst : std_logic := '0';
  signal pd_deb : std_logic;
   constant clk_period : time := 40 ns;
BEGIN
 -- Instantiate VHDL code for button debouncing
   uut: debouncer2 PORT MAP (
          pbutton => pbutton,
          clk => clk,
--          rst => rst,
          pd_deb => pd_deb
        );
   clk_process :process
   begin
  clk <= '0';
  wait for clk_period;
  clk <= '1';
  wait for clk_period;
   end process;
   -- Stimulus process
   stim_proc: process
   begin  
      -- hold reset state for 100 ns.
      wait for 10 ns; 
--      rst <= '1';
      wait for 10 ns; 
--      rst <= '0';
      wait for 100 ns; 

      wait for clk_period*10;
  pbutton <= '0';
  wait for 10 ns; 
  pbutton <= '1';
  wait for 20 ns; 
  pbutton <= '0';
  wait for 10 ns; 
  pbutton <= '1';
  wait for 30 ns; 
  pbutton <= '0';
  wait for 10 ns; 
  pbutton <= '1';
  wait for 40 ns; 
  pbutton <= '0';
  wait for 10 ns; 
  pbutton <= '1';
  wait for 30 ns;  
  pbutton <= '0';
  wait for 10 ns; 
  pbutton <= '1';
  wait for 400 ns;  
  pbutton <= '0';
  wait for 10 ns; 
  pbutton <= '1';
  wait for 20 ns; 
  pbutton <= '0';
  wait for 10 ns; 
  pbutton <= '1';
  wait for 30 ns; 
  pbutton <= '0';
      wait;
   end process;

END;
