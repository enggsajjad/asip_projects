-- VHDL Preprocessor version 0.57
-- module     : 32-bit 3-port multiplexor
-- feature    : select one input from n input ports.
-- references : start from scratch
-- author     : Tak. Tokihisa
-- version    : 1.0  : first cut 2002/01/15
-- VHDL       : 87

-- Functionality : synthesis level
--  port
--   data_in  : input data
--   data_out : selected data 
--   select     : data_out <= data_in0 when sel = "00" else
--            : data_in1 when sel = "01" else
--            : data_in2;



library ieee;
  use ieee.std_logic_1164.all;
  use ieee.std_logic_unsigned.all;
  use ieee.std_logic_arith.all;

entity fhm_multiplexor_w32_00 is
  port (
        data_in0 : in std_logic_vector(31 downto 0);
        data_in1 : in std_logic_vector(31 downto 0);
        data_in2 : in std_logic_vector(31 downto 0);
        sel      : in std_logic_vector(1 downto 0);
        data_out : out std_logic_vector(31 downto 0));
end fhm_multiplexor_w32_00;

architecture synthesis of fhm_multiplexor_w32_00 is
begin
  data_out <= data_in0 when sel = "00" else
	      data_in1 when sel = "01" else
	      data_in2;
end synthesis;

-----------------------------------------
-- Generated by ASIP Meister ver.1.1 --
-----------------------------------------

-----------------------------------------
-- Generated by ASIP Meister ver.1.1 --
-----------------------------------------
