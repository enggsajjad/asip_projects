-----------------------------------------------------------
-- Entity Name: rtg_mux2to1_w1
-----------------------------------------------------------

library IEEE;
use IEEE.std_logic_1164.all;

entity rtg_mux2to1_w1 is
  port (
    SEL : in std_logic;
    DIN0 : in std_logic;
    DIN1 : in std_logic;
    DOUT : out std_logic
  );
end entity rtg_mux2to1_w1;

architecture RTL of rtg_mux2to1_w1 is


begin
  DOUT <= DIN0 when SEL = '0' else 
	DIN1 when SEL = '1' else 
	'X';
end RTL;

-----------------------------------------
-- Generated by ASIP Meister ver.1.1 --
-----------------------------------------

-----------------------------------------
-- Generated by ASIP Meister ver.1.1 --
-----------------------------------------
