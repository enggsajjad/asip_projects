-- Module     : Shifter
-- Feature    : Shift Right or Left, Arithmetic or Logic
-- References : Started from scratch.
-- Author     : Designed by T.Morifuji (c)1996.

-- Version    : 1.1  : Modified by K.Ueda 2001/12/12
--                     Add rotate function
--            : 1.2  : Modified by Y.Yamane 2001/12/26
--            : 1.3  : Modified by Y.Yamane 2001/01/15

-- Comment :
--  mode
--   00  : shift left  logic
--   01  : shift left  arithmetic
--   10  : shift right logic
--   11  : shift right arithmetic

--  ctrl : shift amount


library IEEE;
  use IEEE.std_logic_1164.all;
  use IEEE.std_logic_arith.all;
  use IEEE.std_logic_unsigned.all;

entity fhm_shifter_w32 is
  port (data_in   : in  std_logic_vector(31 downto 0);
        mode      : in  std_logic_vector(1 downto 0);
        ctrl      : in  std_logic_vector(4 downto 0);
        data_out  : out std_logic_vector(31 downto 0));
end fhm_shifter_w32;

architecture synthesis of fhm_shifter_w32 is
  signal int1       : std_logic_vector(31 downto 0);
  signal int2       : std_logic_vector(31 downto 0);
  signal int4       : std_logic_vector(31 downto 0);
  signal int8       : std_logic_vector(31 downto 0);
  signal int16      : std_logic_vector(31 downto 0);
  signal sign1      : std_logic;
  signal sign2      : std_logic_vector(1 downto 0);
  signal sign4      : std_logic_vector(3 downto 0);
  signal sign8      : std_logic_vector(7 downto 0);
  signal sign16     : std_logic_vector(15 downto 0);
  signal rl    : std_logic;
  signal al    : std_logic;
  signal s_cnt : std_logic_vector(4 downto 0);

begin

  s_cnt <= ctrl;
  rl <= mode(1);
  al <= mode(0);

  --  generate sign vectors
  sign1 <= data_in(31) when (al = '1') else
           '0';
  sign2 <= data_in(31) & data_in(31) when (al = '1') else
           (others => '0');
  sign4 <= (3 downto 0 => data_in(31)) when (al = '1') else
           (others => '0');
  sign8 <= (7 downto 0 => data_in(31)) when (al = '1') else
           (others => '0');
  sign16<= (15 downto 0 => data_in(31)) when (al = '1') else
           (others => '0');

  -- 1 bit shift
  first_step: block
  begin  --  block first_step
    int1 <= data_in(30 downto 0) & '0'
			when (s_cnt(0)='1') and (rl = '0') and (al = '0') else
            data_in(31) & data_in(29 downto 0) & '0'
			when (s_cnt(0)='1') and (rl = '0') and (al = '1') else
            sign1 & data_in(31 downto 1) 
			when (s_cnt(0)='1') and (rl = '1') else
            data_in;
  end block first_step;

  -- 2 bit shift
  second_step: block
  begin  --  block second_step 
    int2 <= int1(29 downto 0) & "00"  
			when (s_cnt(1)='1') and (rl = '0') and (al = '0') else
            int1(31) & int1(28 downto 0) & "00"  
			when (s_cnt(1)='1') and (rl = '0') and (al = '1') else
            sign2 & int1(31 downto 2) 
			when (s_cnt(1)='1') and (rl = '1') else
            int1;
  end block second_step;

  -- 4 bit shift
  third_step: block
  begin  --  block third_step 
    int4 <= int2(27 downto 0) & "0000"
			when (s_cnt(2)='1') and (rl = '0') and (al = '0') else
            int2(31) & int2(26 downto 0) & "0000"
			when (s_cnt(2)='1') and (rl = '0') and (al = '1') else
            sign4 & int2(31 downto 4)
			when (s_cnt(2)='1') and (rl = '1') else
            int2;
  end block third_step;

  -- 8 bit shift
  fourth_step: block
  begin  --  block fourth_step 
    int8 <= int4(23 downto 0) & "00000000"
			 when (s_cnt(3)='1') and (rl = '0') and (al = '0') else
            int4(31) & int4(22 downto 0) & "00000000"
			 when (s_cnt(3)='1') and (rl = '0') and (al = '1') else
            sign8 & int4(31 downto 8) 
			 when (s_cnt(3)='1') and (rl = '1') else
            int4;
  end block fourth_step;

  -- 16 bit shift
  fifth_step: block
  begin  --  block fifth_step 
    int16 <= int8(15 downto 0) & "0000000000000000" 
		        when (s_cnt(4)='1') and (rl = '0') and (al = '0') else
             int8(31) & int8(14 downto 0) & "0000000000000000" 
		        when (s_cnt(4)='1') and (rl = '0') and (al = '1') else
             sign16 & int8(31 downto 16) 
		        when (s_cnt(4)='1') and (rl = '1') else
             int8;
  end block fifth_step;

  data_out <= int16;
end synthesis;

-----------------------------------------
-- Generated by ASIP Meister ver.1.1 --
-----------------------------------------
