-- Module     : 1-bit full adder
-- References :
-- Author     : Designed by T.Morifuji (c)1996.
-- Version    : 1.0  :
-- VHDL       : 87

-- Functionality : synthesis level
--  port
--   a, b   : add datas
--   cin    : carry in
--   result : result of a + b + c
--   cout   : carry of a + b + c

library IEEE;
  use IEEE.std_logic_1164.all;
  use IEEE.std_logic_unsigned.all;

entity fhm_adder_w32_fa is
    port (a, b:   in  std_logic;
          cin:    in  std_logic;
          result: out std_logic;
          cout:   out std_logic );
end fhm_adder_w32_fa;

architecture synthesis of fhm_adder_w32_fa is
begin

   result <= (not a and b and not cin) or
	     (a and not b and not cin) or
             (not a and not b and cin) or 
	     (a and b and cin);

   cout <= (a and b and not cin) or 
           (not a and b and cin) or 
           (a and not b and cin) or 
           (a and b and cin);

end synthesis;

--%%

-- Module     : 32-bit ripple carry adder
-- References :
-- Author     : Designed by T.Morifuji (c)1996.
-- Version    : 1.0
-- VHDL       : 87

-- Functionality : synthesis level
--  port
--   a, b   : add datas
--   cin    : carry in
--   result : result of a + b + c
--   cout   : '1' when result > 2^32-1 else '0'

library IEEE;
  use IEEE.std_logic_1164.all;
  use IEEE.std_logic_unsigned.all;

entity fhm_adder_w32 is
    port (a, b   : in  std_logic_vector(31 downto 0);
          cin    : in  std_logic;
          result : out std_logic_vector(31 downto 0);
          cout   : out std_logic);
end fhm_adder_w32;

architecture synthesis of fhm_adder_w32 is

   component fhm_adder_w32_fa
      port (a:      in  std_logic;
            b:      in  std_logic;
            cin:    in  std_logic;
            result: out std_logic;
            cout:   out std_logic);
   end component;

   signal  ctmp :  std_logic_vector(32 downto 0);

begin

   ctmp(0) <= cin;

   full_adder: for i in 31 downto 0 generate
   fan: fhm_adder_w32_fa 
      port map (a      => a(i),
                b      => b(i),
                cin    => ctmp(i),
                result => result(i),
                cout   => ctmp(i+1));
   end generate full_adder;

   cout <= ctmp(32);

end synthesis;

-----------------------------------------
-- Generated by ASIP Meister ver.1.1 --
-----------------------------------------
