-- Module	 : Instruction Memory Access Unit
-- Author	 : M. Itoh (c) 2000.
--                 Modified by K.Ueda (c) 2002
-- Version	 : 1.0
-- VHDL          : 87

-- Functionality : synthesis level
--  port
--    addr     : address from cpu
--    addr_bus : address output for bus
--    data_bus : data from bus
--    data     : data for cpu

library ieee;
use ieee.std_logic_1164.all;

entity fhm_imau_w32 is
  port(
    addr     : in  std_logic_vector(31 downto 0);
    addr_bus : out std_logic_vector(31 downto 0);
    data_bus : in  std_logic_vector(31 downto 0);
    data     : out std_logic_vector(31 downto 0)
  );
end fhm_imau_w32;

architecture synthesis of fhm_imau_w32 is
begin
  addr_bus <= addr;
  data     <= data_bus;
end synthesis;

-----------------------------------------
-- Generated by ASIP Meister ver.1.1 --
-----------------------------------------
