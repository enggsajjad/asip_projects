-- VHDL       : '87
-- Module     : Sign Extender
-- Feature    : extend sign
-- References : Started from scratch.
-- Author     : Tak. Tokihisa
-- Version : 1.0  : 2002/01/14

-- Functionality : synthesis level
--  port
--   data_in  : data extended
--   data_out : extended data 
--   mode     : 0  zero extention
--            : 1  sign extention

library IEEE;
  use IEEE.std_logic_1164.all;
  use IEEE.std_logic_unsigned.all;

entity fhm_extender_w28 is
  port (data_in  : in std_logic_vector(27 downto 0);
        mode     : in std_logic;
        data_out : out std_logic_vector(31 downto 0));
end fhm_extender_w28;

architecture synthesis of fhm_extender_w28 is
begin
  data_out(27 downto 0) <= data_in(27 downto 0);
  sign_ext : for i in 31 downto 28 generate
     data_out(i) <= data_in(27) when mode = '1' else '0';
  end generate sign_ext;
end synthesis;

-----------------------------------------
-- Generated by ASIP Meister ver.1.1 --
-----------------------------------------
